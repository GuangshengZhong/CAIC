`include "src/defines.v"
module Forward_Unit_Id(
    input reg_write_mem,rd_mem,
    input rs1_id,rs2_id,
    input branch_id, jal_id, jalr_id,
    output rs1_fwd_id,rs2_fwd_id
)
endmodule