`include "src/defines.v"
module Forward_Unit_Ex(
    input reg_write_mem,rd_mem,
    input rs1_ex,rs2_ex,
    input reg_write_wb,rd_wb,
    output rs1_fwd_ex,rs2_fwd_ex
)
endmodule
